library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity e_modulo_counter is
	generic( n: natural := 4 );
	port (	sl_clock, sl_reset_n:	in		std_logic;
			sl_enable:				in		std_logic;
			slv_rollover_value:		in		std_logic_vector(n-1 downto 0);
			slv_Q:					out		std_logic_vector(n-1 downto 0);
			sl_rollover:			out		std_logic
	);
end entity e_modulo_counter;

architecture a_modulo_counter of e_modulo_counter is

-- Declarations:

-- Signal Declarations:
	signal u_rollover_value_int:	unsigned(n-1 downto 0):= (others => '0');
	signal u_counter_int:			unsigned(n-1 downto 0):= (others => '0');

begin

-- Assignments:

-- Concurrent Assignments:
	slv_Q <= std_logic_vector(u_counter_int);
	
	u_rollover_value_int <= unsigned(slv_rollover_value);
	
-- Conditional Signal Assignments:
	sl_rollover <= '1' when (u_counter_int = (u_rollover_value_int-1)) else '0';

-- Sequential process with async. low-active reset:
	p_mod_cnt: process(sl_clock, sl_reset_n)
	begin
		if(sl_reset_n = '0') then
			u_counter_int <= (others => '0');
		elsif(rising_edge(sl_clock)) then
			if(sl_enable = '1') then
				if(u_counter_int >= (u_rollover_value_int-1)) then
					u_counter_int <= (others => '0');
				else
					u_counter_int <= u_counter_int + 1;
				end if;
			end if;
		end if;
	end process p_mod_cnt;

end architecture a_modulo_counter;
	